interface adder_intf(input logic clk);
  logic [2:0] a;
  logic [2:0] b;
  logic [3:0] sum;
  logic rst;
endinterface